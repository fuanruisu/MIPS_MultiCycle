module proof();
reg [7:0] mema [0:255];

endmodule 